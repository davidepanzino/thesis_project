/opt/pdk/tsmc28/SRAM/macros/tsdn28hpcpuhdb64x64m4mwa_170a/LEF/tsdn28hpcpuhdb64x64m4mwa_170a.lef