/opt/pdk/tsmc28/SRAM/macros/tsdn28hpcpuhdb64x128m4mwa_170a/LEF/tsdn28hpcpuhdb64x128m4mwa_170a.lef