/opt/pdk/tsmc28/iolib/tpbn28v_160a_FE/TSMCHOME/digital/Back_End/lef/tpbn28v_160a/cup/9m/9M_5X1Y1Z1U/lef/tpbn28v_9lm.lef