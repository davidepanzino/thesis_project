/opt/pdk/tsmc28/SRAM/macros/ts6n28hpcphvta16x16m2fwbso_200b/LEF/ts6n28hpcphvta16x16m2fwbso_200b.lef